
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hd2de7cac;
    ram_cell[       1] = 32'h0;  // 32'h30aaa1ea;
    ram_cell[       2] = 32'h0;  // 32'h6655f6b7;
    ram_cell[       3] = 32'h0;  // 32'h70224917;
    ram_cell[       4] = 32'h0;  // 32'h678c55ec;
    ram_cell[       5] = 32'h0;  // 32'hd40d418e;
    ram_cell[       6] = 32'h0;  // 32'h59593ce5;
    ram_cell[       7] = 32'h0;  // 32'hab564f3c;
    ram_cell[       8] = 32'h0;  // 32'h2b4a21cc;
    ram_cell[       9] = 32'h0;  // 32'h232d7d98;
    ram_cell[      10] = 32'h0;  // 32'hd0194190;
    ram_cell[      11] = 32'h0;  // 32'h4ae6e03b;
    ram_cell[      12] = 32'h0;  // 32'h8c5da8a6;
    ram_cell[      13] = 32'h0;  // 32'hb94041a0;
    ram_cell[      14] = 32'h0;  // 32'hadfac478;
    ram_cell[      15] = 32'h0;  // 32'hdd95a879;
    ram_cell[      16] = 32'h0;  // 32'hf9f3490c;
    ram_cell[      17] = 32'h0;  // 32'hc3fccd41;
    ram_cell[      18] = 32'h0;  // 32'h54a35f8f;
    ram_cell[      19] = 32'h0;  // 32'h2a7f50e0;
    ram_cell[      20] = 32'h0;  // 32'hba7b7dac;
    ram_cell[      21] = 32'h0;  // 32'hec2fb562;
    ram_cell[      22] = 32'h0;  // 32'h9f03e1db;
    ram_cell[      23] = 32'h0;  // 32'h23c658b7;
    ram_cell[      24] = 32'h0;  // 32'h458e447d;
    ram_cell[      25] = 32'h0;  // 32'h9abbdc5e;
    ram_cell[      26] = 32'h0;  // 32'hd07f2bd9;
    ram_cell[      27] = 32'h0;  // 32'h1e963a4f;
    ram_cell[      28] = 32'h0;  // 32'hfbee3003;
    ram_cell[      29] = 32'h0;  // 32'h42b336d2;
    ram_cell[      30] = 32'h0;  // 32'h6500cabe;
    ram_cell[      31] = 32'h0;  // 32'hbc0d6eed;
    ram_cell[      32] = 32'h0;  // 32'h02635574;
    ram_cell[      33] = 32'h0;  // 32'hb40dbc36;
    ram_cell[      34] = 32'h0;  // 32'hb743ee8d;
    ram_cell[      35] = 32'h0;  // 32'h49efd3fd;
    ram_cell[      36] = 32'h0;  // 32'ha4dacfd0;
    ram_cell[      37] = 32'h0;  // 32'h03e23914;
    ram_cell[      38] = 32'h0;  // 32'h483db17d;
    ram_cell[      39] = 32'h0;  // 32'h273f0756;
    ram_cell[      40] = 32'h0;  // 32'hf39941cb;
    ram_cell[      41] = 32'h0;  // 32'h8f925be1;
    ram_cell[      42] = 32'h0;  // 32'hcbfa8c45;
    ram_cell[      43] = 32'h0;  // 32'h81ae44ae;
    ram_cell[      44] = 32'h0;  // 32'h85ca0b91;
    ram_cell[      45] = 32'h0;  // 32'hc32c5d39;
    ram_cell[      46] = 32'h0;  // 32'haaaf2382;
    ram_cell[      47] = 32'h0;  // 32'hac59653e;
    ram_cell[      48] = 32'h0;  // 32'h97552588;
    ram_cell[      49] = 32'h0;  // 32'h0deb1c52;
    ram_cell[      50] = 32'h0;  // 32'hbcb35ab8;
    ram_cell[      51] = 32'h0;  // 32'he319a533;
    ram_cell[      52] = 32'h0;  // 32'h27679a5b;
    ram_cell[      53] = 32'h0;  // 32'ha9e9da72;
    ram_cell[      54] = 32'h0;  // 32'hb86e4e98;
    ram_cell[      55] = 32'h0;  // 32'hd687739f;
    ram_cell[      56] = 32'h0;  // 32'h76f1cfe1;
    ram_cell[      57] = 32'h0;  // 32'hec551743;
    ram_cell[      58] = 32'h0;  // 32'h8b3371f5;
    ram_cell[      59] = 32'h0;  // 32'h91891a59;
    ram_cell[      60] = 32'h0;  // 32'h5e0d17e4;
    ram_cell[      61] = 32'h0;  // 32'h60133b80;
    ram_cell[      62] = 32'h0;  // 32'h09a7f46a;
    ram_cell[      63] = 32'h0;  // 32'h0fe06de9;
    ram_cell[      64] = 32'h0;  // 32'hcf1e4734;
    ram_cell[      65] = 32'h0;  // 32'hf7d5811a;
    ram_cell[      66] = 32'h0;  // 32'h1a33c24a;
    ram_cell[      67] = 32'h0;  // 32'h16584cf8;
    ram_cell[      68] = 32'h0;  // 32'h5d7a64ba;
    ram_cell[      69] = 32'h0;  // 32'h8a2134ea;
    ram_cell[      70] = 32'h0;  // 32'h048e1c72;
    ram_cell[      71] = 32'h0;  // 32'h4cf3b755;
    ram_cell[      72] = 32'h0;  // 32'hb3c141f9;
    ram_cell[      73] = 32'h0;  // 32'h873a7705;
    ram_cell[      74] = 32'h0;  // 32'h43c87844;
    ram_cell[      75] = 32'h0;  // 32'h73ac4a5c;
    ram_cell[      76] = 32'h0;  // 32'h01ea32c4;
    ram_cell[      77] = 32'h0;  // 32'h16347aaf;
    ram_cell[      78] = 32'h0;  // 32'h306178bb;
    ram_cell[      79] = 32'h0;  // 32'h0cafe028;
    ram_cell[      80] = 32'h0;  // 32'h296234f8;
    ram_cell[      81] = 32'h0;  // 32'h1fa3e73f;
    ram_cell[      82] = 32'h0;  // 32'hf03dc65f;
    ram_cell[      83] = 32'h0;  // 32'hcf90aa11;
    ram_cell[      84] = 32'h0;  // 32'h3cb84e3f;
    ram_cell[      85] = 32'h0;  // 32'h16da617a;
    ram_cell[      86] = 32'h0;  // 32'h8c64f717;
    ram_cell[      87] = 32'h0;  // 32'h808f2165;
    ram_cell[      88] = 32'h0;  // 32'h40c4a6cd;
    ram_cell[      89] = 32'h0;  // 32'h421417d3;
    ram_cell[      90] = 32'h0;  // 32'h69c3510b;
    ram_cell[      91] = 32'h0;  // 32'hdc1f9faa;
    ram_cell[      92] = 32'h0;  // 32'hc97995cb;
    ram_cell[      93] = 32'h0;  // 32'h6a68c851;
    ram_cell[      94] = 32'h0;  // 32'h3d38ea8e;
    ram_cell[      95] = 32'h0;  // 32'h025f7d0e;
    ram_cell[      96] = 32'h0;  // 32'h983d9ef4;
    ram_cell[      97] = 32'h0;  // 32'h9b226602;
    ram_cell[      98] = 32'h0;  // 32'h2f49cebd;
    ram_cell[      99] = 32'h0;  // 32'hcf6147f9;
    ram_cell[     100] = 32'h0;  // 32'h066b9680;
    ram_cell[     101] = 32'h0;  // 32'h1640282a;
    ram_cell[     102] = 32'h0;  // 32'hb9787488;
    ram_cell[     103] = 32'h0;  // 32'h6cd3b272;
    ram_cell[     104] = 32'h0;  // 32'h0b5b71fb;
    ram_cell[     105] = 32'h0;  // 32'h848ff03c;
    ram_cell[     106] = 32'h0;  // 32'hd0b5a75e;
    ram_cell[     107] = 32'h0;  // 32'hb9d45cd1;
    ram_cell[     108] = 32'h0;  // 32'h7c5d6937;
    ram_cell[     109] = 32'h0;  // 32'h59e6db2f;
    ram_cell[     110] = 32'h0;  // 32'h3ba24d37;
    ram_cell[     111] = 32'h0;  // 32'h90083e5a;
    ram_cell[     112] = 32'h0;  // 32'hcf094c45;
    ram_cell[     113] = 32'h0;  // 32'h43133c20;
    ram_cell[     114] = 32'h0;  // 32'hb2debd4d;
    ram_cell[     115] = 32'h0;  // 32'h3ecf8f0c;
    ram_cell[     116] = 32'h0;  // 32'hb9cad39c;
    ram_cell[     117] = 32'h0;  // 32'h6a536cd8;
    ram_cell[     118] = 32'h0;  // 32'h4c97e7a5;
    ram_cell[     119] = 32'h0;  // 32'hd5468d4c;
    ram_cell[     120] = 32'h0;  // 32'h78b07af8;
    ram_cell[     121] = 32'h0;  // 32'h7f12f21e;
    ram_cell[     122] = 32'h0;  // 32'h0bb0c139;
    ram_cell[     123] = 32'h0;  // 32'h1c173099;
    ram_cell[     124] = 32'h0;  // 32'hff92b48e;
    ram_cell[     125] = 32'h0;  // 32'h94d4272d;
    ram_cell[     126] = 32'h0;  // 32'hbd81bed5;
    ram_cell[     127] = 32'h0;  // 32'h64b5e9b2;
    ram_cell[     128] = 32'h0;  // 32'h14ed92c5;
    ram_cell[     129] = 32'h0;  // 32'h10747d0d;
    ram_cell[     130] = 32'h0;  // 32'hcca0ea7b;
    ram_cell[     131] = 32'h0;  // 32'hb048a1e6;
    ram_cell[     132] = 32'h0;  // 32'h4ec78ac4;
    ram_cell[     133] = 32'h0;  // 32'h96ee8732;
    ram_cell[     134] = 32'h0;  // 32'h48e6279b;
    ram_cell[     135] = 32'h0;  // 32'h9f4c458a;
    ram_cell[     136] = 32'h0;  // 32'h0fafeadc;
    ram_cell[     137] = 32'h0;  // 32'h9572c044;
    ram_cell[     138] = 32'h0;  // 32'hac7113ec;
    ram_cell[     139] = 32'h0;  // 32'h9b1c041c;
    ram_cell[     140] = 32'h0;  // 32'h9baeb795;
    ram_cell[     141] = 32'h0;  // 32'hdb8ba6d8;
    ram_cell[     142] = 32'h0;  // 32'h8a792576;
    ram_cell[     143] = 32'h0;  // 32'hda6b5022;
    ram_cell[     144] = 32'h0;  // 32'h51c7a24e;
    ram_cell[     145] = 32'h0;  // 32'h945b28ba;
    ram_cell[     146] = 32'h0;  // 32'h8a36c980;
    ram_cell[     147] = 32'h0;  // 32'hf98149e3;
    ram_cell[     148] = 32'h0;  // 32'hf1587c08;
    ram_cell[     149] = 32'h0;  // 32'hdefa9d59;
    ram_cell[     150] = 32'h0;  // 32'h1c969229;
    ram_cell[     151] = 32'h0;  // 32'h0fc3680d;
    ram_cell[     152] = 32'h0;  // 32'hdd6ad658;
    ram_cell[     153] = 32'h0;  // 32'hccffa45c;
    ram_cell[     154] = 32'h0;  // 32'h05c8907f;
    ram_cell[     155] = 32'h0;  // 32'h78355f5f;
    ram_cell[     156] = 32'h0;  // 32'h6bfada93;
    ram_cell[     157] = 32'h0;  // 32'hdca3cc1f;
    ram_cell[     158] = 32'h0;  // 32'h13372cf0;
    ram_cell[     159] = 32'h0;  // 32'hd0462c19;
    ram_cell[     160] = 32'h0;  // 32'h77dc1aa5;
    ram_cell[     161] = 32'h0;  // 32'ha8060482;
    ram_cell[     162] = 32'h0;  // 32'h1a15a592;
    ram_cell[     163] = 32'h0;  // 32'h7276fecd;
    ram_cell[     164] = 32'h0;  // 32'h62551a39;
    ram_cell[     165] = 32'h0;  // 32'h75224527;
    ram_cell[     166] = 32'h0;  // 32'h91155ef4;
    ram_cell[     167] = 32'h0;  // 32'h05cc927c;
    ram_cell[     168] = 32'h0;  // 32'h26a9b281;
    ram_cell[     169] = 32'h0;  // 32'h170e3fcc;
    ram_cell[     170] = 32'h0;  // 32'hd8d5dc3c;
    ram_cell[     171] = 32'h0;  // 32'hbd1a141d;
    ram_cell[     172] = 32'h0;  // 32'h2ccd6d18;
    ram_cell[     173] = 32'h0;  // 32'h04bb08b9;
    ram_cell[     174] = 32'h0;  // 32'hf76d0473;
    ram_cell[     175] = 32'h0;  // 32'h20696089;
    ram_cell[     176] = 32'h0;  // 32'hba50f385;
    ram_cell[     177] = 32'h0;  // 32'he6fd37ea;
    ram_cell[     178] = 32'h0;  // 32'h4df721f1;
    ram_cell[     179] = 32'h0;  // 32'h7e46f613;
    ram_cell[     180] = 32'h0;  // 32'hcac3c50c;
    ram_cell[     181] = 32'h0;  // 32'h53b54bd2;
    ram_cell[     182] = 32'h0;  // 32'haadbdb7b;
    ram_cell[     183] = 32'h0;  // 32'h4065e27f;
    ram_cell[     184] = 32'h0;  // 32'h4e7ebde4;
    ram_cell[     185] = 32'h0;  // 32'h1b306aea;
    ram_cell[     186] = 32'h0;  // 32'h386e4793;
    ram_cell[     187] = 32'h0;  // 32'h7e9893af;
    ram_cell[     188] = 32'h0;  // 32'hf2a9470a;
    ram_cell[     189] = 32'h0;  // 32'h013a840f;
    ram_cell[     190] = 32'h0;  // 32'h9efd41ae;
    ram_cell[     191] = 32'h0;  // 32'hcf3fd009;
    ram_cell[     192] = 32'h0;  // 32'h46d42b40;
    ram_cell[     193] = 32'h0;  // 32'he3983e8f;
    ram_cell[     194] = 32'h0;  // 32'hb29cbdff;
    ram_cell[     195] = 32'h0;  // 32'hcd6552e7;
    ram_cell[     196] = 32'h0;  // 32'h3789b3de;
    ram_cell[     197] = 32'h0;  // 32'h4be66654;
    ram_cell[     198] = 32'h0;  // 32'h18c89bde;
    ram_cell[     199] = 32'h0;  // 32'h6ebe9130;
    ram_cell[     200] = 32'h0;  // 32'ha373e1ad;
    ram_cell[     201] = 32'h0;  // 32'h8e7b2192;
    ram_cell[     202] = 32'h0;  // 32'h0ef83d5c;
    ram_cell[     203] = 32'h0;  // 32'h65520b82;
    ram_cell[     204] = 32'h0;  // 32'h0a926b35;
    ram_cell[     205] = 32'h0;  // 32'ha9a590b6;
    ram_cell[     206] = 32'h0;  // 32'h04655828;
    ram_cell[     207] = 32'h0;  // 32'h584412a0;
    ram_cell[     208] = 32'h0;  // 32'h07653688;
    ram_cell[     209] = 32'h0;  // 32'h6e7f25f5;
    ram_cell[     210] = 32'h0;  // 32'h9ca70513;
    ram_cell[     211] = 32'h0;  // 32'h0c1fa118;
    ram_cell[     212] = 32'h0;  // 32'heb1028bf;
    ram_cell[     213] = 32'h0;  // 32'h333d91a3;
    ram_cell[     214] = 32'h0;  // 32'hff0b4039;
    ram_cell[     215] = 32'h0;  // 32'h6089d41c;
    ram_cell[     216] = 32'h0;  // 32'h35031827;
    ram_cell[     217] = 32'h0;  // 32'h43999b38;
    ram_cell[     218] = 32'h0;  // 32'h8508cdb2;
    ram_cell[     219] = 32'h0;  // 32'h5302d2a9;
    ram_cell[     220] = 32'h0;  // 32'hbdda1b04;
    ram_cell[     221] = 32'h0;  // 32'h24340ccb;
    ram_cell[     222] = 32'h0;  // 32'h4e7ddafd;
    ram_cell[     223] = 32'h0;  // 32'h230a5314;
    ram_cell[     224] = 32'h0;  // 32'h118d458f;
    ram_cell[     225] = 32'h0;  // 32'h860c7a7b;
    ram_cell[     226] = 32'h0;  // 32'hd370e669;
    ram_cell[     227] = 32'h0;  // 32'h1070ff9c;
    ram_cell[     228] = 32'h0;  // 32'he3fea50f;
    ram_cell[     229] = 32'h0;  // 32'h1b903dc9;
    ram_cell[     230] = 32'h0;  // 32'h947e5956;
    ram_cell[     231] = 32'h0;  // 32'h8251a87c;
    ram_cell[     232] = 32'h0;  // 32'h95f56c04;
    ram_cell[     233] = 32'h0;  // 32'hb0204feb;
    ram_cell[     234] = 32'h0;  // 32'h046eb424;
    ram_cell[     235] = 32'h0;  // 32'he23b11ad;
    ram_cell[     236] = 32'h0;  // 32'he565a19f;
    ram_cell[     237] = 32'h0;  // 32'h639ef331;
    ram_cell[     238] = 32'h0;  // 32'h2a8962e5;
    ram_cell[     239] = 32'h0;  // 32'h3cadf555;
    ram_cell[     240] = 32'h0;  // 32'h6d120137;
    ram_cell[     241] = 32'h0;  // 32'h135e8726;
    ram_cell[     242] = 32'h0;  // 32'h35e5f2a7;
    ram_cell[     243] = 32'h0;  // 32'ha6d56371;
    ram_cell[     244] = 32'h0;  // 32'h6a18c078;
    ram_cell[     245] = 32'h0;  // 32'h06582b0f;
    ram_cell[     246] = 32'h0;  // 32'haa29acdc;
    ram_cell[     247] = 32'h0;  // 32'hb2b0e516;
    ram_cell[     248] = 32'h0;  // 32'hd506887a;
    ram_cell[     249] = 32'h0;  // 32'hd94787ae;
    ram_cell[     250] = 32'h0;  // 32'hec7a61f5;
    ram_cell[     251] = 32'h0;  // 32'h062c793a;
    ram_cell[     252] = 32'h0;  // 32'h6aab6124;
    ram_cell[     253] = 32'h0;  // 32'h1dd8f61f;
    ram_cell[     254] = 32'h0;  // 32'hfe1a888d;
    ram_cell[     255] = 32'h0;  // 32'h41ed2d75;
    // src matrix A
    ram_cell[     256] = 32'h05b94784;
    ram_cell[     257] = 32'h331036f2;
    ram_cell[     258] = 32'he67ddfe6;
    ram_cell[     259] = 32'h317476c5;
    ram_cell[     260] = 32'ha1370d9c;
    ram_cell[     261] = 32'h20e945bc;
    ram_cell[     262] = 32'h4f8d392e;
    ram_cell[     263] = 32'hef8df8ca;
    ram_cell[     264] = 32'h10d62861;
    ram_cell[     265] = 32'hc0a491c8;
    ram_cell[     266] = 32'hdbdaf493;
    ram_cell[     267] = 32'ha3225fa3;
    ram_cell[     268] = 32'h9171579d;
    ram_cell[     269] = 32'h3487c579;
    ram_cell[     270] = 32'h02393eed;
    ram_cell[     271] = 32'h131d5cec;
    ram_cell[     272] = 32'h3a700656;
    ram_cell[     273] = 32'he669d0ae;
    ram_cell[     274] = 32'hb352ddaf;
    ram_cell[     275] = 32'hcce498f0;
    ram_cell[     276] = 32'h1c4d8199;
    ram_cell[     277] = 32'hdf84ebf5;
    ram_cell[     278] = 32'h3e002f8c;
    ram_cell[     279] = 32'he507fc75;
    ram_cell[     280] = 32'h4b61c81a;
    ram_cell[     281] = 32'h75c07fd6;
    ram_cell[     282] = 32'h71a5387d;
    ram_cell[     283] = 32'h79a83331;
    ram_cell[     284] = 32'hf2a70ea7;
    ram_cell[     285] = 32'h9bbf9a20;
    ram_cell[     286] = 32'hffaffee5;
    ram_cell[     287] = 32'hf1dc521d;
    ram_cell[     288] = 32'h6f613ab6;
    ram_cell[     289] = 32'h3524f46f;
    ram_cell[     290] = 32'h9c8d1ac2;
    ram_cell[     291] = 32'hb0c90edf;
    ram_cell[     292] = 32'h2564c8b2;
    ram_cell[     293] = 32'h61f2021f;
    ram_cell[     294] = 32'h7e3c0358;
    ram_cell[     295] = 32'h0c9fac7f;
    ram_cell[     296] = 32'h43a212f2;
    ram_cell[     297] = 32'h68cb6eb5;
    ram_cell[     298] = 32'h63e58258;
    ram_cell[     299] = 32'he76d328e;
    ram_cell[     300] = 32'he1725c71;
    ram_cell[     301] = 32'he136e492;
    ram_cell[     302] = 32'h901c6c16;
    ram_cell[     303] = 32'h3b40a66f;
    ram_cell[     304] = 32'h4a9222bb;
    ram_cell[     305] = 32'h64c3fac6;
    ram_cell[     306] = 32'hfdf5d3a3;
    ram_cell[     307] = 32'hd10912ab;
    ram_cell[     308] = 32'h86febd0d;
    ram_cell[     309] = 32'h7d20a9fd;
    ram_cell[     310] = 32'hb40f8e8f;
    ram_cell[     311] = 32'haf6b8714;
    ram_cell[     312] = 32'h1620fabe;
    ram_cell[     313] = 32'h34594f77;
    ram_cell[     314] = 32'h8c8b4717;
    ram_cell[     315] = 32'h5e05e0f1;
    ram_cell[     316] = 32'h77f6fdb3;
    ram_cell[     317] = 32'h61a95232;
    ram_cell[     318] = 32'hff113e5b;
    ram_cell[     319] = 32'ha9000720;
    ram_cell[     320] = 32'h2649d57a;
    ram_cell[     321] = 32'h687152f1;
    ram_cell[     322] = 32'hb5757650;
    ram_cell[     323] = 32'h35c6a39c;
    ram_cell[     324] = 32'h122f936c;
    ram_cell[     325] = 32'h4a80fad1;
    ram_cell[     326] = 32'hf7921910;
    ram_cell[     327] = 32'h6266112b;
    ram_cell[     328] = 32'hecf9d9bc;
    ram_cell[     329] = 32'hcc32afcb;
    ram_cell[     330] = 32'hcd598bec;
    ram_cell[     331] = 32'hdc8310f7;
    ram_cell[     332] = 32'h125d2032;
    ram_cell[     333] = 32'hfc1a75ac;
    ram_cell[     334] = 32'hf4d90b0a;
    ram_cell[     335] = 32'h220d4fda;
    ram_cell[     336] = 32'h6c5fb01c;
    ram_cell[     337] = 32'hce67f43c;
    ram_cell[     338] = 32'h920dd390;
    ram_cell[     339] = 32'ha6d98efd;
    ram_cell[     340] = 32'h6c08d268;
    ram_cell[     341] = 32'h15146780;
    ram_cell[     342] = 32'hecdeda4e;
    ram_cell[     343] = 32'ha370da2e;
    ram_cell[     344] = 32'h986f8cc1;
    ram_cell[     345] = 32'h5d98a3a0;
    ram_cell[     346] = 32'ha23becaa;
    ram_cell[     347] = 32'hf369c58a;
    ram_cell[     348] = 32'he8f05766;
    ram_cell[     349] = 32'h609ef128;
    ram_cell[     350] = 32'hef28e5fc;
    ram_cell[     351] = 32'h0906fdf2;
    ram_cell[     352] = 32'h16d4f73f;
    ram_cell[     353] = 32'h8968c07a;
    ram_cell[     354] = 32'h44b935a5;
    ram_cell[     355] = 32'h14774bfc;
    ram_cell[     356] = 32'h21421ddf;
    ram_cell[     357] = 32'h0adf7822;
    ram_cell[     358] = 32'hc727b9a9;
    ram_cell[     359] = 32'h87a94d85;
    ram_cell[     360] = 32'hdfc75e57;
    ram_cell[     361] = 32'h727eaf6a;
    ram_cell[     362] = 32'h2a04cf9d;
    ram_cell[     363] = 32'h967e0051;
    ram_cell[     364] = 32'h0ca5d80a;
    ram_cell[     365] = 32'h9e035842;
    ram_cell[     366] = 32'h62da30d7;
    ram_cell[     367] = 32'h3b639658;
    ram_cell[     368] = 32'h9f44bcf1;
    ram_cell[     369] = 32'h00a70100;
    ram_cell[     370] = 32'h3d972b89;
    ram_cell[     371] = 32'h1f443f89;
    ram_cell[     372] = 32'h43536e5f;
    ram_cell[     373] = 32'he9eae332;
    ram_cell[     374] = 32'h935821ed;
    ram_cell[     375] = 32'h6fdc645c;
    ram_cell[     376] = 32'he300296f;
    ram_cell[     377] = 32'h7562401e;
    ram_cell[     378] = 32'h9bc7907e;
    ram_cell[     379] = 32'hd5fe82a5;
    ram_cell[     380] = 32'ha3c68d0e;
    ram_cell[     381] = 32'ha050f642;
    ram_cell[     382] = 32'he8346267;
    ram_cell[     383] = 32'hd847e5a5;
    ram_cell[     384] = 32'h4d2c2e67;
    ram_cell[     385] = 32'h38a4156e;
    ram_cell[     386] = 32'hc8a17c9e;
    ram_cell[     387] = 32'h729cba09;
    ram_cell[     388] = 32'heea9eaee;
    ram_cell[     389] = 32'hfe4a32af;
    ram_cell[     390] = 32'h15f97769;
    ram_cell[     391] = 32'hfe931aa5;
    ram_cell[     392] = 32'heb966452;
    ram_cell[     393] = 32'h60edb076;
    ram_cell[     394] = 32'hf2d43769;
    ram_cell[     395] = 32'ha0a8f252;
    ram_cell[     396] = 32'h8a862a78;
    ram_cell[     397] = 32'h32f964e9;
    ram_cell[     398] = 32'h33753163;
    ram_cell[     399] = 32'hbebb49ed;
    ram_cell[     400] = 32'he7b214e1;
    ram_cell[     401] = 32'h96c9ad1b;
    ram_cell[     402] = 32'h16301727;
    ram_cell[     403] = 32'h8996a032;
    ram_cell[     404] = 32'h6786940f;
    ram_cell[     405] = 32'h092729a8;
    ram_cell[     406] = 32'h525af7a8;
    ram_cell[     407] = 32'hf11b46c6;
    ram_cell[     408] = 32'hb2819418;
    ram_cell[     409] = 32'h0481e9ef;
    ram_cell[     410] = 32'hfca2d9b9;
    ram_cell[     411] = 32'hc832f820;
    ram_cell[     412] = 32'h055e09e2;
    ram_cell[     413] = 32'h4f61bbde;
    ram_cell[     414] = 32'h9ea69f1c;
    ram_cell[     415] = 32'h3831e0fc;
    ram_cell[     416] = 32'he58d89ae;
    ram_cell[     417] = 32'h3a150b60;
    ram_cell[     418] = 32'h399cacf9;
    ram_cell[     419] = 32'h5aaef7d2;
    ram_cell[     420] = 32'h01982230;
    ram_cell[     421] = 32'hcab78376;
    ram_cell[     422] = 32'h68c7deab;
    ram_cell[     423] = 32'hea96bafe;
    ram_cell[     424] = 32'h632752f8;
    ram_cell[     425] = 32'haceec87a;
    ram_cell[     426] = 32'h05192d0b;
    ram_cell[     427] = 32'he4ee24e8;
    ram_cell[     428] = 32'he4c8fda6;
    ram_cell[     429] = 32'h73f4f9e9;
    ram_cell[     430] = 32'heeb67e9d;
    ram_cell[     431] = 32'h31a766d5;
    ram_cell[     432] = 32'h9dc5da79;
    ram_cell[     433] = 32'h1d334ec7;
    ram_cell[     434] = 32'hbf561cd1;
    ram_cell[     435] = 32'h47ee8063;
    ram_cell[     436] = 32'h15ce3b31;
    ram_cell[     437] = 32'h18ba3901;
    ram_cell[     438] = 32'habb23139;
    ram_cell[     439] = 32'hc76df968;
    ram_cell[     440] = 32'h05aad2f6;
    ram_cell[     441] = 32'h998169c3;
    ram_cell[     442] = 32'hde530867;
    ram_cell[     443] = 32'heeae1b8f;
    ram_cell[     444] = 32'h99f66500;
    ram_cell[     445] = 32'h23bd06e6;
    ram_cell[     446] = 32'h58f9b5fb;
    ram_cell[     447] = 32'h5a37c442;
    ram_cell[     448] = 32'h17841eb3;
    ram_cell[     449] = 32'h225cdc6e;
    ram_cell[     450] = 32'ha6ba575e;
    ram_cell[     451] = 32'h1f005f9f;
    ram_cell[     452] = 32'h191320fa;
    ram_cell[     453] = 32'hf8131b95;
    ram_cell[     454] = 32'h348a47fe;
    ram_cell[     455] = 32'hf2ca04cf;
    ram_cell[     456] = 32'hd29651fb;
    ram_cell[     457] = 32'hde0ce7bc;
    ram_cell[     458] = 32'h84a3537a;
    ram_cell[     459] = 32'h0de95491;
    ram_cell[     460] = 32'hf23424bd;
    ram_cell[     461] = 32'he65f1a3b;
    ram_cell[     462] = 32'h41dd9963;
    ram_cell[     463] = 32'hce0d12f2;
    ram_cell[     464] = 32'h5854b46c;
    ram_cell[     465] = 32'hc62fe223;
    ram_cell[     466] = 32'hf704ae1e;
    ram_cell[     467] = 32'h4ff77537;
    ram_cell[     468] = 32'h49e037d9;
    ram_cell[     469] = 32'h5e2f14e3;
    ram_cell[     470] = 32'hb7fe10e7;
    ram_cell[     471] = 32'h6fa448b9;
    ram_cell[     472] = 32'hfc16d085;
    ram_cell[     473] = 32'hab86ac82;
    ram_cell[     474] = 32'hc594e07b;
    ram_cell[     475] = 32'hd86b6b56;
    ram_cell[     476] = 32'h8da7af21;
    ram_cell[     477] = 32'h990e85e2;
    ram_cell[     478] = 32'hc45c502c;
    ram_cell[     479] = 32'h7ac1a449;
    ram_cell[     480] = 32'hab8ef5ef;
    ram_cell[     481] = 32'hba1bd912;
    ram_cell[     482] = 32'h1a5bcd39;
    ram_cell[     483] = 32'h96027517;
    ram_cell[     484] = 32'hd4831024;
    ram_cell[     485] = 32'hd828c26f;
    ram_cell[     486] = 32'h68fd65c6;
    ram_cell[     487] = 32'h6dc0fb7b;
    ram_cell[     488] = 32'h8c795b14;
    ram_cell[     489] = 32'hea6172f4;
    ram_cell[     490] = 32'h10495dd0;
    ram_cell[     491] = 32'h29b3841c;
    ram_cell[     492] = 32'h4eacbb46;
    ram_cell[     493] = 32'h00aad771;
    ram_cell[     494] = 32'h4cbb1abb;
    ram_cell[     495] = 32'h433a282a;
    ram_cell[     496] = 32'h1c93a583;
    ram_cell[     497] = 32'h563657bf;
    ram_cell[     498] = 32'he2f805c0;
    ram_cell[     499] = 32'hf17c55ba;
    ram_cell[     500] = 32'h7662e36d;
    ram_cell[     501] = 32'h4e5c75d3;
    ram_cell[     502] = 32'h04ea97bb;
    ram_cell[     503] = 32'h8ba4a13f;
    ram_cell[     504] = 32'h7f5d53db;
    ram_cell[     505] = 32'h4a0c6649;
    ram_cell[     506] = 32'h9e2596a2;
    ram_cell[     507] = 32'h47324100;
    ram_cell[     508] = 32'he66b0675;
    ram_cell[     509] = 32'h787350c4;
    ram_cell[     510] = 32'hebe8bcb8;
    ram_cell[     511] = 32'h2ea36574;
    // src matrix B
    ram_cell[     512] = 32'h1375b9b3;
    ram_cell[     513] = 32'hf07609cc;
    ram_cell[     514] = 32'hc8235cdd;
    ram_cell[     515] = 32'h31da5ebb;
    ram_cell[     516] = 32'hc4198c50;
    ram_cell[     517] = 32'h3aefd55f;
    ram_cell[     518] = 32'hf05851d7;
    ram_cell[     519] = 32'h78c7068a;
    ram_cell[     520] = 32'hf1e2d0b0;
    ram_cell[     521] = 32'heb211e0d;
    ram_cell[     522] = 32'h3fcfc4b4;
    ram_cell[     523] = 32'he1d0a5c8;
    ram_cell[     524] = 32'h35a11a13;
    ram_cell[     525] = 32'hc8d632f9;
    ram_cell[     526] = 32'h9c91b403;
    ram_cell[     527] = 32'hcd5523fe;
    ram_cell[     528] = 32'h9b00f682;
    ram_cell[     529] = 32'h5b0c23ff;
    ram_cell[     530] = 32'h9a03c09b;
    ram_cell[     531] = 32'h51c25ae0;
    ram_cell[     532] = 32'hf277810e;
    ram_cell[     533] = 32'h73fdcbca;
    ram_cell[     534] = 32'hc360391e;
    ram_cell[     535] = 32'hb4a4f69c;
    ram_cell[     536] = 32'h7f46d2c7;
    ram_cell[     537] = 32'h45e0e68e;
    ram_cell[     538] = 32'hc27af355;
    ram_cell[     539] = 32'h3b58cc78;
    ram_cell[     540] = 32'h36338eec;
    ram_cell[     541] = 32'h80b9bb2d;
    ram_cell[     542] = 32'h80127a84;
    ram_cell[     543] = 32'hdf22bbc3;
    ram_cell[     544] = 32'hb0706725;
    ram_cell[     545] = 32'h63fa34a3;
    ram_cell[     546] = 32'h5f177533;
    ram_cell[     547] = 32'h17bbe439;
    ram_cell[     548] = 32'hdaa2ffb8;
    ram_cell[     549] = 32'heb29a55a;
    ram_cell[     550] = 32'haabe4431;
    ram_cell[     551] = 32'h06889843;
    ram_cell[     552] = 32'h4b2b58ba;
    ram_cell[     553] = 32'h942e6432;
    ram_cell[     554] = 32'h5a32b6e8;
    ram_cell[     555] = 32'h91066220;
    ram_cell[     556] = 32'h804fd692;
    ram_cell[     557] = 32'hca95fd56;
    ram_cell[     558] = 32'hd1e60835;
    ram_cell[     559] = 32'h25202599;
    ram_cell[     560] = 32'hefbed348;
    ram_cell[     561] = 32'h512ba33c;
    ram_cell[     562] = 32'hd9674ba9;
    ram_cell[     563] = 32'hc854ce10;
    ram_cell[     564] = 32'h3be4c744;
    ram_cell[     565] = 32'h055f56e9;
    ram_cell[     566] = 32'h31c3e77f;
    ram_cell[     567] = 32'h1c9383a9;
    ram_cell[     568] = 32'hd9590e27;
    ram_cell[     569] = 32'h4dbc0e7b;
    ram_cell[     570] = 32'h44bb6af0;
    ram_cell[     571] = 32'h432d0fbf;
    ram_cell[     572] = 32'hb5436367;
    ram_cell[     573] = 32'hf53c22c4;
    ram_cell[     574] = 32'h585265da;
    ram_cell[     575] = 32'h66a781f8;
    ram_cell[     576] = 32'he1f1be6e;
    ram_cell[     577] = 32'ha8a7d42f;
    ram_cell[     578] = 32'ha0ac015a;
    ram_cell[     579] = 32'h521bef83;
    ram_cell[     580] = 32'h2bcd03ad;
    ram_cell[     581] = 32'h3dd1cc3d;
    ram_cell[     582] = 32'hcabba163;
    ram_cell[     583] = 32'h3374a11e;
    ram_cell[     584] = 32'hcbf21dd5;
    ram_cell[     585] = 32'h074f785d;
    ram_cell[     586] = 32'ha879a733;
    ram_cell[     587] = 32'h37cff90e;
    ram_cell[     588] = 32'hdf6c71a8;
    ram_cell[     589] = 32'he4bd2e0c;
    ram_cell[     590] = 32'h999438d6;
    ram_cell[     591] = 32'hba7084c6;
    ram_cell[     592] = 32'h234adfca;
    ram_cell[     593] = 32'h964a8529;
    ram_cell[     594] = 32'hc9b14979;
    ram_cell[     595] = 32'ha13b8e5e;
    ram_cell[     596] = 32'h042a94e2;
    ram_cell[     597] = 32'he128cb25;
    ram_cell[     598] = 32'he7ce4769;
    ram_cell[     599] = 32'h43f907c4;
    ram_cell[     600] = 32'hca07022b;
    ram_cell[     601] = 32'hf931a430;
    ram_cell[     602] = 32'h9824b44b;
    ram_cell[     603] = 32'h42fdc2c3;
    ram_cell[     604] = 32'h75c11e64;
    ram_cell[     605] = 32'h4b6271f1;
    ram_cell[     606] = 32'h25f8105a;
    ram_cell[     607] = 32'hbea65851;
    ram_cell[     608] = 32'h1f7b61d0;
    ram_cell[     609] = 32'hb1c40882;
    ram_cell[     610] = 32'h5d73c535;
    ram_cell[     611] = 32'h56c513bb;
    ram_cell[     612] = 32'h17eb8a56;
    ram_cell[     613] = 32'h25fb8d3c;
    ram_cell[     614] = 32'he944b1df;
    ram_cell[     615] = 32'hfdd39b9a;
    ram_cell[     616] = 32'haf943573;
    ram_cell[     617] = 32'h8d962884;
    ram_cell[     618] = 32'h74717356;
    ram_cell[     619] = 32'h28d6d61f;
    ram_cell[     620] = 32'h94d5afa7;
    ram_cell[     621] = 32'h657031ec;
    ram_cell[     622] = 32'h91af934b;
    ram_cell[     623] = 32'h7760b02b;
    ram_cell[     624] = 32'hf9096282;
    ram_cell[     625] = 32'h344d2f17;
    ram_cell[     626] = 32'h805c385f;
    ram_cell[     627] = 32'hcc58e1a1;
    ram_cell[     628] = 32'he9f1997d;
    ram_cell[     629] = 32'h2c1afc1c;
    ram_cell[     630] = 32'h93f40545;
    ram_cell[     631] = 32'hfb0af3d6;
    ram_cell[     632] = 32'he699ee6d;
    ram_cell[     633] = 32'h8199fd88;
    ram_cell[     634] = 32'h9437be09;
    ram_cell[     635] = 32'hc4f23973;
    ram_cell[     636] = 32'h7cd747e3;
    ram_cell[     637] = 32'h1771d23d;
    ram_cell[     638] = 32'h47a461d1;
    ram_cell[     639] = 32'h747c67e7;
    ram_cell[     640] = 32'hb46079ce;
    ram_cell[     641] = 32'hb5f9fd15;
    ram_cell[     642] = 32'h3d136280;
    ram_cell[     643] = 32'hc7631811;
    ram_cell[     644] = 32'h2ee36b0f;
    ram_cell[     645] = 32'hdbe1bfdb;
    ram_cell[     646] = 32'hee3777b2;
    ram_cell[     647] = 32'h296a3ae2;
    ram_cell[     648] = 32'h7b2d1750;
    ram_cell[     649] = 32'hbe921c0a;
    ram_cell[     650] = 32'hb7c7f71f;
    ram_cell[     651] = 32'h4b19a397;
    ram_cell[     652] = 32'h2f2c886e;
    ram_cell[     653] = 32'hec91d2ef;
    ram_cell[     654] = 32'h2c579eae;
    ram_cell[     655] = 32'h22229bb6;
    ram_cell[     656] = 32'hbc03b6c5;
    ram_cell[     657] = 32'h4eb0f412;
    ram_cell[     658] = 32'hd796d73c;
    ram_cell[     659] = 32'h4a478ffe;
    ram_cell[     660] = 32'h82b47840;
    ram_cell[     661] = 32'he8578ab5;
    ram_cell[     662] = 32'h73279760;
    ram_cell[     663] = 32'hf8cb7efa;
    ram_cell[     664] = 32'hbf101c43;
    ram_cell[     665] = 32'h2d93c7f5;
    ram_cell[     666] = 32'h3e084f8f;
    ram_cell[     667] = 32'hd344885a;
    ram_cell[     668] = 32'haf2acaef;
    ram_cell[     669] = 32'h2e76276e;
    ram_cell[     670] = 32'hb1a49b74;
    ram_cell[     671] = 32'h0055c564;
    ram_cell[     672] = 32'hf81e9b9b;
    ram_cell[     673] = 32'hcb2cd793;
    ram_cell[     674] = 32'haa675fff;
    ram_cell[     675] = 32'h34a4f40e;
    ram_cell[     676] = 32'h015ad5f9;
    ram_cell[     677] = 32'h51670494;
    ram_cell[     678] = 32'h30daad3c;
    ram_cell[     679] = 32'hb6c57702;
    ram_cell[     680] = 32'ha8182211;
    ram_cell[     681] = 32'h61efcf71;
    ram_cell[     682] = 32'h7217cb40;
    ram_cell[     683] = 32'h80d412f5;
    ram_cell[     684] = 32'h696a516f;
    ram_cell[     685] = 32'hc61ebb05;
    ram_cell[     686] = 32'h975ddd34;
    ram_cell[     687] = 32'hb142b4ab;
    ram_cell[     688] = 32'h678596ab;
    ram_cell[     689] = 32'h85fc0059;
    ram_cell[     690] = 32'h9db57933;
    ram_cell[     691] = 32'h409c8531;
    ram_cell[     692] = 32'hd6546207;
    ram_cell[     693] = 32'hc1ce5966;
    ram_cell[     694] = 32'he64db8f2;
    ram_cell[     695] = 32'he5af9123;
    ram_cell[     696] = 32'hd5a977cf;
    ram_cell[     697] = 32'hc8a43924;
    ram_cell[     698] = 32'he902a3ca;
    ram_cell[     699] = 32'h76fac9ee;
    ram_cell[     700] = 32'h75d5a982;
    ram_cell[     701] = 32'h5f27ed26;
    ram_cell[     702] = 32'h27167894;
    ram_cell[     703] = 32'h1cdf94e5;
    ram_cell[     704] = 32'h83840567;
    ram_cell[     705] = 32'h17f4d499;
    ram_cell[     706] = 32'hfeb4ee60;
    ram_cell[     707] = 32'hb0a38490;
    ram_cell[     708] = 32'h494b21f3;
    ram_cell[     709] = 32'h8a6bcf6e;
    ram_cell[     710] = 32'h54ee713b;
    ram_cell[     711] = 32'h30679614;
    ram_cell[     712] = 32'h8e204712;
    ram_cell[     713] = 32'h094e5085;
    ram_cell[     714] = 32'h4ce8d831;
    ram_cell[     715] = 32'h139141e2;
    ram_cell[     716] = 32'h97b2f754;
    ram_cell[     717] = 32'h74109338;
    ram_cell[     718] = 32'h820f308e;
    ram_cell[     719] = 32'ha910f79d;
    ram_cell[     720] = 32'h775162c3;
    ram_cell[     721] = 32'hb7aacd04;
    ram_cell[     722] = 32'h11e5d115;
    ram_cell[     723] = 32'hf0137815;
    ram_cell[     724] = 32'hea9c18b7;
    ram_cell[     725] = 32'h94d85905;
    ram_cell[     726] = 32'hdaa5abb2;
    ram_cell[     727] = 32'h4b5e7fb8;
    ram_cell[     728] = 32'h40e83293;
    ram_cell[     729] = 32'h8641f95a;
    ram_cell[     730] = 32'h1fdfbf95;
    ram_cell[     731] = 32'h21005fa5;
    ram_cell[     732] = 32'h17a5b165;
    ram_cell[     733] = 32'h80e36909;
    ram_cell[     734] = 32'h7d6e92dd;
    ram_cell[     735] = 32'h027b9f6d;
    ram_cell[     736] = 32'hc998268e;
    ram_cell[     737] = 32'h6c3de7f2;
    ram_cell[     738] = 32'h1cfa242f;
    ram_cell[     739] = 32'hacad46d6;
    ram_cell[     740] = 32'h325a68f9;
    ram_cell[     741] = 32'h81522c37;
    ram_cell[     742] = 32'hb8fd99bf;
    ram_cell[     743] = 32'h9f49c1a0;
    ram_cell[     744] = 32'h1a4b25a8;
    ram_cell[     745] = 32'h57eba163;
    ram_cell[     746] = 32'h56c2cdcb;
    ram_cell[     747] = 32'hb68ba61b;
    ram_cell[     748] = 32'h4d85ad29;
    ram_cell[     749] = 32'he53be63f;
    ram_cell[     750] = 32'hf9b14ae9;
    ram_cell[     751] = 32'ha7860a15;
    ram_cell[     752] = 32'h836a2d38;
    ram_cell[     753] = 32'h68fc6398;
    ram_cell[     754] = 32'hde413645;
    ram_cell[     755] = 32'h975db610;
    ram_cell[     756] = 32'heb482e1c;
    ram_cell[     757] = 32'hbed014ad;
    ram_cell[     758] = 32'had6c706d;
    ram_cell[     759] = 32'hef80cdd5;
    ram_cell[     760] = 32'h74e9f6e2;
    ram_cell[     761] = 32'h3def43ba;
    ram_cell[     762] = 32'h6be61912;
    ram_cell[     763] = 32'hf088f4b5;
    ram_cell[     764] = 32'hc0cb9232;
    ram_cell[     765] = 32'h22e166fe;
    ram_cell[     766] = 32'h8a69e5e3;
    ram_cell[     767] = 32'ha1867cf4;
end

endmodule

